module Top(
    input   i_clk,
    input   i_rst_n
);

 
parameter T         =   50;
parameter fg        =   1;
parameter fs        =   0.5;
parameter fc        =   1;
parameter maxLen    =   16;
parameter minLen    =   4;
parameter brushR    =   {4'd8, 4'd4, 4'd2};


endmodule